module progmem (
    // Closk & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,
    input  wire [31:0] addr,
    output wire [31:0] rdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 10;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin

  mem['h0000] <= 32'h20010737;
  mem['h0001] <= 32'h02030537;
  mem['h0002] <= 32'h010008b7;
  mem['h0003] <= 32'haaaab5b7;
  mem['h0004] <= 32'h00002637;
  mem['h0005] <= 32'h10350513;
  mem['h0006] <= 32'h00000793;
  mem['h0007] <= 32'hffa88893;
  mem['h0008] <= 32'h00780337;
  mem['h0009] <= 32'h01c70813;
  mem['h000A] <= 32'haaa58593;
  mem['h000B] <= 32'h71060613;
  mem['h000C] <= 32'h0180006f;
  mem['h000D] <= 32'h00672223;
  mem['h000E] <= 32'h00b82023;
  mem['h000F] <= 32'h00a72023;
  mem['h0010] <= 32'h00178793;
  mem['h0011] <= 32'h02c78063;
  mem['h0012] <= 32'h0017f693;
  mem['h0013] <= 32'hfe0684e3;
  mem['h0014] <= 32'h01172223;
  mem['h0015] <= 32'h00b82023;
  mem['h0016] <= 32'h00a72023;
  mem['h0017] <= 32'h00178793;
  mem['h0018] <= 32'hfec794e3;
  mem['h0019] <= 32'h0000006f;
  mem['h001A] <= 32'h200007b7;
  mem['h001B] <= 32'h0047a503;
  mem['h001C] <= 32'h00157513;
  mem['h001D] <= 32'h00008067;
  mem['h001E] <= 32'h20000737;
  mem['h001F] <= 32'h00472783;
  mem['h0020] <= 32'h0017f793;
  mem['h0021] <= 32'hfe079ce3;
  mem['h0022] <= 32'h00a72623;
  mem['h0023] <= 32'h00008067;
  mem['h0024] <= 32'h00054683;
  mem['h0025] <= 32'h02068263;
  mem['h0026] <= 32'h20000737;
  mem['h0027] <= 32'h00150513;
  mem['h0028] <= 32'h00472783;
  mem['h0029] <= 32'h0017f793;
  mem['h002A] <= 32'hfe079ce3;
  mem['h002B] <= 32'h00d72623;
  mem['h002C] <= 32'h00054683;
  mem['h002D] <= 32'hfe0694e3;
  mem['h002E] <= 32'h00008067;
  mem['h002F] <= 32'hfc010113;
  mem['h0030] <= 32'h00054303;
  mem['h0031] <= 32'h02f12a23;
  mem['h0032] <= 32'h02410793;
  mem['h0033] <= 32'h02b12223;
  mem['h0034] <= 32'h02c12423;
  mem['h0035] <= 32'h02d12623;
  mem['h0036] <= 32'h02e12823;
  mem['h0037] <= 32'h03012c23;
  mem['h0038] <= 32'h03112e23;
  mem['h0039] <= 32'h00f12423;
  mem['h003A] <= 32'h06030a63;
  mem['h003B] <= 32'h00150613;
  mem['h003C] <= 32'h00000693;
  mem['h003D] <= 32'h00000e13;
  mem['h003E] <= 32'h00000793;
  mem['h003F] <= 32'h02500593;
  mem['h0040] <= 32'h20000737;
  mem['h0041] <= 32'h00a00893;
  mem['h0042] <= 32'h04800813;
  mem['h0043] <= 32'h00000517;
  mem['h0044] <= 32'h44850513;
  mem['h0045] <= 32'h04078863;
  mem['h0046] <= 32'hfd030313;
  mem['h0047] <= 32'h0ff37313;
  mem['h0048] <= 32'h00686c63;
  mem['h0049] <= 32'h00231313;
  mem['h004A] <= 32'h00a30333;
  mem['h004B] <= 32'h00032303;
  mem['h004C] <= 32'h00a30333;
  mem['h004D] <= 32'h00030067;
  mem['h004E] <= 32'h00472783;
  mem['h004F] <= 32'h0017f793;
  mem['h0050] <= 32'hfe079ce3;
  mem['h0051] <= 32'h00b72623;
  mem['h0052] <= 32'h00000693;
  mem['h0053] <= 32'h00000e13;
  mem['h0054] <= 32'h00064303;
  mem['h0055] <= 32'h00160613;
  mem['h0056] <= 32'hfa031ee3;
  mem['h0057] <= 32'h04010113;
  mem['h0058] <= 32'h00008067;
  mem['h0059] <= 32'h00100793;
  mem['h005A] <= 32'hfeb304e3;
  mem['h005B] <= 32'h00472783;
  mem['h005C] <= 32'h0017f793;
  mem['h005D] <= 32'hfe079ce3;
  mem['h005E] <= 32'h00672623;
  mem['h005F] <= 32'hfd131ae3;
  mem['h0060] <= 32'h20000337;
  mem['h0061] <= 32'h00432783;
  mem['h0062] <= 32'h0017f793;
  mem['h0063] <= 32'hfe079ce3;
  mem['h0064] <= 32'h00d00e93;
  mem['h0065] <= 32'h01d32623;
  mem['h0066] <= 32'hfb9ff06f;
  mem['h0067] <= 32'h00812783;
  mem['h0068] <= 32'h00478e93;
  mem['h0069] <= 32'h1e0e0263;
  mem['h006A] <= 32'h0007a283;
  mem['h006B] <= 32'h01d12423;
  mem['h006C] <= 32'h01c00313;
  mem['h006D] <= 32'h00900f93;
  mem['h006E] <= 32'h200006b7;
  mem['h006F] <= 32'hffc00f13;
  mem['h0070] <= 32'h0062d7b3;
  mem['h0071] <= 32'h00f7fe93;
  mem['h0072] <= 32'h057e8e13;
  mem['h0073] <= 32'h01dfe463;
  mem['h0074] <= 32'h030e8e13;
  mem['h0075] <= 32'h0046a783;
  mem['h0076] <= 32'h0017f793;
  mem['h0077] <= 32'hfe079ce3;
  mem['h0078] <= 32'h01c6a623;
  mem['h0079] <= 32'hffc30313;
  mem['h007A] <= 32'hfde31ce3;
  mem['h007B] <= 32'h00000693;
  mem['h007C] <= 32'h00000e13;
  mem['h007D] <= 32'h00000793;
  mem['h007E] <= 32'hf59ff06f;
  mem['h007F] <= 32'h00812783;
  mem['h0080] <= 32'h0007a303;
  mem['h0081] <= 32'h00478793;
  mem['h0082] <= 32'h00f12423;
  mem['h0083] <= 32'h00034e03;
  mem['h0084] <= 32'hfc0e0ee3;
  mem['h0085] <= 32'h200006b7;
  mem['h0086] <= 32'h00130313;
  mem['h0087] <= 32'h0046a783;
  mem['h0088] <= 32'h0017f793;
  mem['h0089] <= 32'hfe079ce3;
  mem['h008A] <= 32'h01c6a623;
  mem['h008B] <= 32'h00034e03;
  mem['h008C] <= 32'hfe0e14e3;
  mem['h008D] <= 32'h00000693;
  mem['h008E] <= 32'h00000e13;
  mem['h008F] <= 32'h00000793;
  mem['h0090] <= 32'hf11ff06f;
  mem['h0091] <= 32'h00812783;
  mem['h0092] <= 32'h00478693;
  mem['h0093] <= 32'h0007a783;
  mem['h0094] <= 32'h00d12423;
  mem['h0095] <= 32'h00a00693;
  mem['h0096] <= 32'h00078e93;
  mem['h0097] <= 32'h02d7c7b3;
  mem['h0098] <= 32'h18078063;
  mem['h0099] <= 32'h00100693;
  mem['h009A] <= 32'h00a00e13;
  mem['h009B] <= 32'h03c7c7b3;
  mem['h009C] <= 32'h00068313;
  mem['h009D] <= 32'h00168693;
  mem['h009E] <= 32'hfe079ae3;
  mem['h009F] <= 32'h00a00f13;
  mem['h00A0] <= 32'h200006b7;
  mem['h00A1] <= 32'hfff00f93;
  mem['h00A2] <= 32'h03eefe33;
  mem['h00A3] <= 32'h030e0e13;
  mem['h00A4] <= 32'h0046a783;
  mem['h00A5] <= 32'h0017f793;
  mem['h00A6] <= 32'hfe079ce3;
  mem['h00A7] <= 32'h01c6a623;
  mem['h00A8] <= 32'hfff30313;
  mem['h00A9] <= 32'h03eedeb3;
  mem['h00AA] <= 32'hfff310e3;
  mem['h00AB] <= 32'h00000693;
  mem['h00AC] <= 32'h00000e13;
  mem['h00AD] <= 32'h00000793;
  mem['h00AE] <= 32'he99ff06f;
  mem['h00AF] <= 32'h00812783;
  mem['h00B0] <= 32'h0007ae03;
  mem['h00B1] <= 32'h00478693;
  mem['h00B2] <= 32'h00d12423;
  mem['h00B3] <= 32'h0e0e4a63;
  mem['h00B4] <= 32'h00a00693;
  mem['h00B5] <= 32'h02de46b3;
  mem['h00B6] <= 32'h10068863;
  mem['h00B7] <= 32'h00100e93;
  mem['h00B8] <= 32'h00a00313;
  mem['h00B9] <= 32'h0266c6b3;
  mem['h00BA] <= 32'h000e8793;
  mem['h00BB] <= 32'h001e8e93;
  mem['h00BC] <= 32'hfe069ae3;
  mem['h00BD] <= 32'h00c10f13;
  mem['h00BE] <= 32'h00ff07b3;
  mem['h00BF] <= 32'h000f0313;
  mem['h00C0] <= 32'h00a00f93;
  mem['h00C1] <= 32'h03fe66b3;
  mem['h00C2] <= 32'h00078293;
  mem['h00C3] <= 32'hfff78793;
  mem['h00C4] <= 32'h03068693;
  mem['h00C5] <= 32'h00d780a3;
  mem['h00C6] <= 32'h03fe4e33;
  mem['h00C7] <= 32'hfe5f14e3;
  mem['h00C8] <= 32'h01df0f33;
  mem['h00C9] <= 32'h200006b7;
  mem['h00CA] <= 32'h00034e03;
  mem['h00CB] <= 32'h0046a783;
  mem['h00CC] <= 32'h0017f793;
  mem['h00CD] <= 32'hfe079ce3;
  mem['h00CE] <= 32'h01c6a623;
  mem['h00CF] <= 32'h00130313;
  mem['h00D0] <= 32'hfe6f14e3;
  mem['h00D1] <= 32'h00000693;
  mem['h00D2] <= 32'h00000e13;
  mem['h00D3] <= 32'h00000793;
  mem['h00D4] <= 32'he01ff06f;
  mem['h00D5] <= 32'h00812783;
  mem['h00D6] <= 32'h200006b7;
  mem['h00D7] <= 32'h0007a303;
  mem['h00D8] <= 32'h00478793;
  mem['h00D9] <= 32'h00f12423;
  mem['h00DA] <= 32'h0046a783;
  mem['h00DB] <= 32'h0017f793;
  mem['h00DC] <= 32'hfe079ce3;
  mem['h00DD] <= 32'h0ff37313;
  mem['h00DE] <= 32'h0066a623;
  mem['h00DF] <= 32'h00000e13;
  mem['h00E0] <= 32'h00000693;
  mem['h00E1] <= 32'hdcdff06f;
  mem['h00E2] <= 32'h00d03333;
  mem['h00E3] <= 32'h40600333;
  mem['h00E4] <= 32'hfe837313;
  mem['h00E5] <= 32'h0007a283;
  mem['h00E6] <= 32'h01d12423;
  mem['h00E7] <= 32'h01c30313;
  mem['h00E8] <= 32'he15ff06f;
  mem['h00E9] <= 32'h00078e13;
  mem['h00EA] <= 32'h00000693;
  mem['h00EB] <= 32'hda5ff06f;
  mem['h00EC] <= 32'h00078693;
  mem['h00ED] <= 32'h00000e13;
  mem['h00EE] <= 32'h00000793;
  mem['h00EF] <= 32'hd95ff06f;
  mem['h00F0] <= 32'h41c00e33;
  mem['h00F1] <= 32'h200006b7;
  mem['h00F2] <= 32'h0046a783;
  mem['h00F3] <= 32'h0017f793;
  mem['h00F4] <= 32'hfe079ce3;
  mem['h00F5] <= 32'h02d00793;
  mem['h00F6] <= 32'h00f6a623;
  mem['h00F7] <= 32'hef5ff06f;
  mem['h00F8] <= 32'h00000313;
  mem['h00F9] <= 32'he99ff06f;
  mem['h00FA] <= 32'h00000793;
  mem['h00FB] <= 32'h00100e93;
  mem['h00FC] <= 32'hf05ff06f;
  mem['h00FD] <= 32'h200007b7;
  mem['h00FE] <= 32'h0047a503;
  mem['h00FF] <= 32'h00355513;
  mem['h0100] <= 32'h00157513;
  mem['h0101] <= 32'h00008067;
  mem['h0102] <= 32'h20000737;
  mem['h0103] <= 32'h00472783;
  mem['h0104] <= 32'h0037d793;
  mem['h0105] <= 32'h0017f793;
  mem['h0106] <= 32'hfe079ae3;
  mem['h0107] <= 32'h00872503;
  mem['h0108] <= 32'h0ff57513;
  mem['h0109] <= 32'h00008067;
  mem['h010A] <= 32'h00050313;
  mem['h010B] <= 32'h20000737;
  mem['h010C] <= 32'h00000513;
  mem['h010D] <= 32'h00800893;
  mem['h010E] <= 32'h00d00e13;
  mem['h010F] <= 32'h05e00e93;
  mem['h0110] <= 32'hfff58f13;
  mem['h0111] <= 32'h00472783;
  mem['h0112] <= 32'h0037d793;
  mem['h0113] <= 32'h0017f793;
  mem['h0114] <= 32'hfe079ae3;
  mem['h0115] <= 32'h00872583;
  mem['h0116] <= 32'h0ff5f693;
  mem['h0117] <= 32'h03168663;
  mem['h0118] <= 32'h03c68e63;
  mem['h0119] <= 32'hfe068793;
  mem['h011A] <= 32'h0ff7f793;
  mem['h011B] <= 32'hfcfeece3;
  mem['h011C] <= 32'hfde55ae3;
  mem['h011D] <= 32'h06061a63;
  mem['h011E] <= 32'h00d30023;
  mem['h011F] <= 32'h00150513;
  mem['h0120] <= 32'h00130313;
  mem['h0121] <= 32'hfc1ff06f;
  mem['h0122] <= 32'hfa050ee3;
  mem['h0123] <= 32'h02061863;
  mem['h0124] <= 32'hfff30313;
  mem['h0125] <= 32'hfff50513;
  mem['h0126] <= 32'hfadff06f;
  mem['h0127] <= 32'h00030023;
  mem['h0128] <= 32'h20000737;
  mem['h0129] <= 32'h00472783;
  mem['h012A] <= 32'h0017f793;
  mem['h012B] <= 32'hfe079ce3;
  mem['h012C] <= 32'h00a00793;
  mem['h012D] <= 32'h00f72623;
  mem['h012E] <= 32'h00008067;
  mem['h012F] <= 32'h00000817;
  mem['h0130] <= 32'h1bc80813;
  mem['h0131] <= 32'h200005b7;
  mem['h0132] <= 32'h00180813;
  mem['h0133] <= 32'h0045a783;
  mem['h0134] <= 32'h0017f793;
  mem['h0135] <= 32'hfe079ce3;
  mem['h0136] <= 32'h00d5a623;
  mem['h0137] <= 32'h00084683;
  mem['h0138] <= 32'hfe0694e3;
  mem['h0139] <= 32'hfadff06f;
  mem['h013A] <= 32'h20000837;
  mem['h013B] <= 32'h00482783;
  mem['h013C] <= 32'h0017f793;
  mem['h013D] <= 32'hfe079ce3;
  mem['h013E] <= 32'h0ff5f593;
  mem['h013F] <= 32'h00b82623;
  mem['h0140] <= 32'hf79ff06f;
  mem['h0141] <= 32'h00054783;
  mem['h0142] <= 32'h00158593;
  mem['h0143] <= 32'h00150513;
  mem['h0144] <= 32'hfff5c703;
  mem['h0145] <= 32'h00078863;
  mem['h0146] <= 32'hfee786e3;
  mem['h0147] <= 32'h40e78533;
  mem['h0148] <= 32'h00008067;
  mem['h0149] <= 32'h40e00533;
  mem['h014A] <= 32'h00008067;
  mem['h014B] <= 32'h00054783;
  mem['h014C] <= 32'h00078e63;
  mem['h014D] <= 32'h00050793;
  mem['h014E] <= 32'h0017c703;
  mem['h014F] <= 32'h00178793;
  mem['h0150] <= 32'hfe071ce3;
  mem['h0151] <= 32'h40a78533;
  mem['h0152] <= 32'h00008067;
  mem['h0153] <= 32'h00000513;
  mem['h0154] <= 32'h00008067;
  mem['h0155] <= 32'hfffffbfc;
  mem['h0156] <= 32'hfffffbfc;
  mem['h0157] <= 32'hfffffbfc;
  mem['h0158] <= 32'hfffffbfc;
  mem['h0159] <= 32'hfffffbfc;
  mem['h015A] <= 32'hfffffbfc;
  mem['h015B] <= 32'hfffffbfc;
  mem['h015C] <= 32'hfffffbfc;
  mem['h015D] <= 32'hfffffbfc;
  mem['h015E] <= 32'hfffffbfc;
  mem['h015F] <= 32'hfffffbe4;
  mem['h0160] <= 32'hfffffbe4;
  mem['h0161] <= 32'hfffffbe4;
  mem['h0162] <= 32'hfffffbe4;
  mem['h0163] <= 32'hfffffbe4;
  mem['h0164] <= 32'hfffffbe4;
  mem['h0165] <= 32'hfffffbe4;
  mem['h0166] <= 32'hfffffbe4;
  mem['h0167] <= 32'hfffffbe4;
  mem['h0168] <= 32'hfffffbe4;
  mem['h0169] <= 32'hfffffbe4;
  mem['h016A] <= 32'hfffffbe4;
  mem['h016B] <= 32'hfffffbe4;
  mem['h016C] <= 32'hfffffbe4;
  mem['h016D] <= 32'hfffffbe4;
  mem['h016E] <= 32'hfffffbe4;
  mem['h016F] <= 32'hfffffbe4;
  mem['h0170] <= 32'hfffffbe4;
  mem['h0171] <= 32'hfffffbe4;
  mem['h0172] <= 32'hfffffbe4;
  mem['h0173] <= 32'hfffffbe4;
  mem['h0174] <= 32'hfffffbe4;
  mem['h0175] <= 32'hfffffbe4;
  mem['h0176] <= 32'hfffffbe4;
  mem['h0177] <= 32'hfffffbe4;
  mem['h0178] <= 32'hfffffbe4;
  mem['h0179] <= 32'hfffffbe4;
  mem['h017A] <= 32'hfffffbe4;
  mem['h017B] <= 32'hfffffbe4;
  mem['h017C] <= 32'hfffffbe4;
  mem['h017D] <= 32'hfffffbe4;
  mem['h017E] <= 32'hfffffbe4;
  mem['h017F] <= 32'hfffffbe4;
  mem['h0180] <= 32'hfffffbe4;
  mem['h0181] <= 32'hfffffbe4;
  mem['h0182] <= 32'hfffffbe4;
  mem['h0183] <= 32'hfffffbe4;
  mem['h0184] <= 32'hfffffbe4;
  mem['h0185] <= 32'hfffffbe4;
  mem['h0186] <= 32'hfffffbe4;
  mem['h0187] <= 32'hfffffbe4;
  mem['h0188] <= 32'hfffffe00;
  mem['h0189] <= 32'hfffffd68;
  mem['h018A] <= 32'hfffffbe4;
  mem['h018B] <= 32'hfffffc48;
  mem['h018C] <= 32'hfffffbe4;
  mem['h018D] <= 32'hfffffe5c;
  mem['h018E] <= 32'hfffffbe4;
  mem['h018F] <= 32'hfffffbe4;
  mem['h0190] <= 32'hfffffbe4;
  mem['h0191] <= 32'hfffffe50;
  mem['h0192] <= 32'hfffffbe4;
  mem['h0193] <= 32'hfffffbe4;
  mem['h0194] <= 32'hfffffbe4;
  mem['h0195] <= 32'hfffffbe4;
  mem['h0196] <= 32'hfffffbe4;
  mem['h0197] <= 32'hfffffbe4;
  mem['h0198] <= 32'hfffffca8;
  mem['h0199] <= 32'hfffffbe4;
  mem['h019A] <= 32'hfffffcf0;
  mem['h019B] <= 32'hfffffbe4;
  mem['h019C] <= 32'hfffffbe4;
  mem['h019D] <= 32'hfffffc48;
  mem['h019E] <= 32'h00082008;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule

