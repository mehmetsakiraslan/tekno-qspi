@40000000
37 07 02 02 B7 07 01 20 13 07 F7 19 23 A0 E7 00
B7 06 01 20 93 07 70 3E 23 A0 E6 00 93 87 F7 FF
E3 9C 07 FE 6F 00 00 00
