@40000000
B7 06 01 20 37 07 04 02 B7 B5 AA AA 13 07 37 10
93 07 00 00 93 08 00 0A 13 88 C6 01 93 85 A5 AA
13 05 80 3E 6F 00 C0 01 23 A2 16 01 23 20 B8 00
23 A0 E6 00 03 A6 86 00 93 87 17 00 63 82 A7 02
13 F6 17 00 E3 02 06 FE 23 A2 06 00 23 20 B8 00
23 A0 E6 00 03 A6 86 00 93 87 17 00 E3 92 A7 FE
B7 07 00 02 93 87 67 10 37 07 01 02 23 A0 F6 00
13 07 57 10 23 A0 E6 00 93 07 30 06 B7 06 01 20
23 A0 E6 00 93 87 F7 FF E3 9C 07 FE B7 B7 AA 1A
93 87 37 AA 23 A4 F6 00 B7 07 00 BC 93 87 F7 FF
23 A6 F6 00 B7 C7 AD DE 93 87 F7 EE 23 A8 F6 00
B7 27 FF FF 93 87 F7 FF 23 AA F6 00 B7 B7 AA 3A
93 87 A7 AA 23 AC F6 00 B7 07 00 60 93 87 77 FF
23 AE F6 00 B7 B7 AA 4A 93 87 67 AA 23 A0 F6 02
B7 A7 E2 24 93 87 57 65 23 A2 F6 02 93 07 00 0B
23 A2 F6 00 B7 07 04 02 93 87 27 50 37 07 01 02
23 A0 F6 00 13 07 57 10 23 A0 E6 00 83 A7 86 00
63 8A 07 00 B7 07 01 20 23 A0 E7 00 83 A6 87 00
E3 9C 06 FE 37 07 01 02 B7 07 01 20 13 07 57 10
23 A0 E7 00 B7 06 01 20 93 07 30 06 23 A0 E6 00
93 87 F7 FF E3 9C 07 FE 37 07 04 02 93 07 00 0D
13 07 37 10 23 A2 F6 00 23 A0 E6 00 6F 00 00 00
B7 07 00 20 03 A5 47 00 13 75 15 00 67 80 00 00
37 07 00 20 83 27 47 00 93 F7 17 00 E3 9C 07 FE
23 26 A7 00 67 80 00 00 83 46 05 00 63 82 06 02
37 07 00 20 13 05 15 00 83 27 47 00 93 F7 17 00
E3 9C 07 FE 23 26 D7 00 83 46 05 00 E3 94 06 FE
67 80 00 00 13 01 01 FC 03 43 05 00 23 2A F1 02
93 07 41 02 23 22 B1 02 23 24 C1 02 23 26 D1 02
23 28 E1 02 23 2C 01 03 23 2E 11 03 23 24 F1 00
63 0A 03 06 13 06 15 00 93 06 00 00 13 0E 00 00
93 07 00 00 93 05 50 02 37 07 00 20 93 08 A0 00
13 08 80 04 17 05 00 00 13 05 85 44 63 88 07 04
13 03 03 FD 13 73 F3 0F 63 6C 68 00 13 13 23 00
33 03 A3 00 03 23 03 00 33 03 A3 00 67 00 03 00
83 27 47 00 93 F7 17 00 E3 9C 07 FE 23 26 B7 00
93 06 00 00 13 0E 00 00 03 43 06 00 13 06 16 00
E3 1E 03 FA 13 01 01 04 67 80 00 00 93 07 10 00
E3 04 B3 FE 83 27 47 00 93 F7 17 00 E3 9C 07 FE
23 26 67 00 E3 1A 13 FD 37 03 00 20 83 27 43 00
93 F7 17 00 E3 9C 07 FE 93 0E D0 00 23 26 D3 01
6F F0 9F FB 83 27 81 00 93 8E 47 00 63 02 0E 1E
83 A2 07 00 23 24 D1 01 13 03 C0 01 93 0F 90 00
B7 06 00 20 13 0F C0 FF B3 D7 62 00 93 FE F7 00
13 8E 7E 05 63 E4 DF 01 13 8E 0E 03 83 A7 46 00
93 F7 17 00 E3 9C 07 FE 23 A6 C6 01 13 03 C3 FF
E3 1C E3 FD 93 06 00 00 13 0E 00 00 93 07 00 00
6F F0 9F F5 83 27 81 00 03 A3 07 00 93 87 47 00
23 24 F1 00 03 4E 03 00 E3 0E 0E FC B7 06 00 20
13 03 13 00 83 A7 46 00 93 F7 17 00 E3 9C 07 FE
23 A6 C6 01 03 4E 03 00 E3 14 0E FE 93 06 00 00
13 0E 00 00 93 07 00 00 6F F0 1F F1 83 27 81 00
93 86 47 00 83 A7 07 00 23 24 D1 00 93 06 A0 00
93 8E 07 00 B3 C7 D7 02 63 80 07 18 93 06 10 00
13 0E A0 00 B3 C7 C7 03 13 83 06 00 93 86 16 00
E3 9A 07 FE 13 0F A0 00 B7 06 00 20 93 0F F0 FF
33 FE EE 03 13 0E 0E 03 83 A7 46 00 93 F7 17 00
E3 9C 07 FE 23 A6 C6 01 13 03 F3 FF B3 DE EE 03
E3 10 F3 FF 93 06 00 00 13 0E 00 00 93 07 00 00
6F F0 9F E9 83 27 81 00 03 AE 07 00 93 86 47 00
23 24 D1 00 63 4A 0E 0E 93 06 A0 00 B3 46 DE 02
63 88 06 10 93 0E 10 00 13 03 A0 00 B3 C6 66 02
93 87 0E 00 93 8E 1E 00 E3 9A 06 FE 13 0F C1 00
B3 07 FF 00 13 03 0F 00 93 0F A0 00 B3 66 FE 03
93 82 07 00 93 87 F7 FF 93 86 06 03 A3 80 D7 00
33 4E FE 03 E3 14 5F FE 33 0F DF 01 B7 06 00 20
03 4E 03 00 83 A7 46 00 93 F7 17 00 E3 9C 07 FE
23 A6 C6 01 13 03 13 00 E3 14 6F FE 93 06 00 00
13 0E 00 00 93 07 00 00 6F F0 1F E0 83 27 81 00
B7 06 00 20 03 A3 07 00 93 87 47 00 23 24 F1 00
83 A7 46 00 93 F7 17 00 E3 9C 07 FE 13 73 F3 0F
23 A6 66 00 13 0E 00 00 93 06 00 00 6F F0 DF DC
33 33 D0 00 33 03 60 40 13 73 83 FE 83 A2 07 00
23 24 D1 01 13 03 C3 01 6F F0 5F E1 13 8E 07 00
93 06 00 00 6F F0 5F DA 93 86 07 00 13 0E 00 00
93 07 00 00 6F F0 5F D9 33 0E C0 41 B7 06 00 20
83 A7 46 00 93 F7 17 00 E3 9C 07 FE 93 07 D0 02
23 A6 F6 00 6F F0 5F EF 13 03 00 00 6F F0 9F E9
93 07 00 00 93 0E 10 00 6F F0 5F F0 B7 07 00 20
03 A5 47 00 13 55 35 00 13 75 15 00 67 80 00 00
37 07 00 20 83 27 47 00 93 D7 37 00 93 F7 17 00
E3 9A 07 FE 03 25 87 00 13 75 F5 0F 67 80 00 00
13 03 05 00 37 07 00 20 13 05 00 00 93 08 80 00
13 0E D0 00 93 0E E0 05 13 8F F5 FF 83 27 47 00
93 D7 37 00 93 F7 17 00 E3 9A 07 FE 83 25 87 00
93 F6 F5 0F 63 86 16 03 63 8E C6 03 93 87 06 FE
93 F7 F7 0F E3 EC FE FC E3 5A E5 FD 63 1A 06 06
23 00 D3 00 13 05 15 00 13 03 13 00 6F F0 1F FC
E3 0E 05 FA 63 18 06 02 13 03 F3 FF 13 05 F5 FF
6F F0 DF FA 23 00 03 00 37 07 00 20 83 27 47 00
93 F7 17 00 E3 9C 07 FE 93 07 A0 00 23 26 F7 00
67 80 00 00 17 08 00 00 13 08 C8 1B B7 05 00 20
13 08 18 00 83 A7 45 00 93 F7 17 00 E3 9C 07 FE
23 A6 D5 00 83 46 08 00 E3 94 06 FE 6F F0 DF FA
37 08 00 20 83 27 48 00 93 F7 17 00 E3 9C 07 FE
93 F5 F5 0F 23 26 B8 00 6F F0 9F F7 83 47 05 00
93 85 15 00 13 05 15 00 03 C7 F5 FF 63 88 07 00
E3 86 E7 FE 33 85 E7 40 67 80 00 00 33 05 E0 40
67 80 00 00 83 47 05 00 63 8E 07 00 93 07 05 00
03 C7 17 00 93 87 17 00 E3 1C 07 FE 33 85 A7 40
67 80 00 00 13 05 00 00 67 80 00 00
@4000064C
FC FB FF FF FC FB FF FF FC FB FF FF FC FB FF FF
FC FB FF FF FC FB FF FF FC FB FF FF FC FB FF FF
FC FB FF FF FC FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF 00 FE FF FF
68 FD FF FF E4 FB FF FF 48 FC FF FF E4 FB FF FF
5C FE FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
50 FE FF FF E4 FB FF FF E4 FB FF FF E4 FB FF FF
E4 FB FF FF E4 FB FF FF E4 FB FF FF A8 FC FF FF
E4 FB FF FF F0 FC FF FF E4 FB FF FF E4 FB FF FF
48 FC FF FF
@40000770
08 20 08 00
