@40000000
B7 B7 AA AA 37 07 01 20 93 87 A7 AA 23 24 F7 00
B7 07 02 02 93 87 F7 19 23 20 F7 00 6F 00 00 00
